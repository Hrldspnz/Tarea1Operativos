// platform.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module platform (
		input  wire       button_external_connection_export,          //          button_external_connection.export
		input  wire       clk_clk,                                    //                                 clk.clk
		output wire [6:0] id7_segmentos_1_external_connection_export, // id7_segmentos_1_external_connection.export
		output wire [6:0] id7_segmentos_2_external_connection_export, // id7_segmentos_2_external_connection.export
		output wire [6:0] id7_segmentos_3_external_connection_export, // id7_segmentos_3_external_connection.export
		output wire [6:0] id7_segmentos_4_external_connection_export, // id7_segmentos_4_external_connection.export
		input  wire       reset_reset_n,                              //                               reset.reset_n
		output wire [6:0] segmentos_5_external_connection_export,     //     segmentos_5_external_connection.export
		output wire [6:0] segmentos_6_external_connection_export,     //     segmentos_6_external_connection.export
		input  wire [1:0] switchs_external_connection_export          //         switchs_external_connection.export
	);

	wire  [31:0] cpu_data_master_readdata;                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [20:0] cpu_data_master_address;                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;         // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;           // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_s1_address;            // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;         // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;              // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;          // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;              // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_segmentos_1_s1_chipselect; // mm_interconnect_0:segmentos_1_s1_chipselect -> segmentos_1:chipselect
	wire  [31:0] mm_interconnect_0_segmentos_1_s1_readdata;   // segmentos_1:readdata -> mm_interconnect_0:segmentos_1_s1_readdata
	wire   [1:0] mm_interconnect_0_segmentos_1_s1_address;    // mm_interconnect_0:segmentos_1_s1_address -> segmentos_1:address
	wire         mm_interconnect_0_segmentos_1_s1_write;      // mm_interconnect_0:segmentos_1_s1_write -> segmentos_1:write_n
	wire  [31:0] mm_interconnect_0_segmentos_1_s1_writedata;  // mm_interconnect_0:segmentos_1_s1_writedata -> segmentos_1:writedata
	wire         mm_interconnect_0_segmentos_2_s1_chipselect; // mm_interconnect_0:segmentos_2_s1_chipselect -> segmentos_2:chipselect
	wire  [31:0] mm_interconnect_0_segmentos_2_s1_readdata;   // segmentos_2:readdata -> mm_interconnect_0:segmentos_2_s1_readdata
	wire   [1:0] mm_interconnect_0_segmentos_2_s1_address;    // mm_interconnect_0:segmentos_2_s1_address -> segmentos_2:address
	wire         mm_interconnect_0_segmentos_2_s1_write;      // mm_interconnect_0:segmentos_2_s1_write -> segmentos_2:write_n
	wire  [31:0] mm_interconnect_0_segmentos_2_s1_writedata;  // mm_interconnect_0:segmentos_2_s1_writedata -> segmentos_2:writedata
	wire         mm_interconnect_0_segmentos_3_s1_chipselect; // mm_interconnect_0:segmentos_3_s1_chipselect -> segmentos_3:chipselect
	wire  [31:0] mm_interconnect_0_segmentos_3_s1_readdata;   // segmentos_3:readdata -> mm_interconnect_0:segmentos_3_s1_readdata
	wire   [1:0] mm_interconnect_0_segmentos_3_s1_address;    // mm_interconnect_0:segmentos_3_s1_address -> segmentos_3:address
	wire         mm_interconnect_0_segmentos_3_s1_write;      // mm_interconnect_0:segmentos_3_s1_write -> segmentos_3:write_n
	wire  [31:0] mm_interconnect_0_segmentos_3_s1_writedata;  // mm_interconnect_0:segmentos_3_s1_writedata -> segmentos_3:writedata
	wire         mm_interconnect_0_segmentos_4_s1_chipselect; // mm_interconnect_0:segmentos_4_s1_chipselect -> segmentos_4:chipselect
	wire  [31:0] mm_interconnect_0_segmentos_4_s1_readdata;   // segmentos_4:readdata -> mm_interconnect_0:segmentos_4_s1_readdata
	wire   [1:0] mm_interconnect_0_segmentos_4_s1_address;    // mm_interconnect_0:segmentos_4_s1_address -> segmentos_4:address
	wire         mm_interconnect_0_segmentos_4_s1_write;      // mm_interconnect_0:segmentos_4_s1_write -> segmentos_4:write_n
	wire  [31:0] mm_interconnect_0_segmentos_4_s1_writedata;  // mm_interconnect_0:segmentos_4_s1_writedata -> segmentos_4:writedata
	wire  [31:0] mm_interconnect_0_switchs_s1_readdata;       // switchs:readdata -> mm_interconnect_0:switchs_s1_readdata
	wire   [1:0] mm_interconnect_0_switchs_s1_address;        // mm_interconnect_0:switchs_s1_address -> switchs:address
	wire         mm_interconnect_0_timer_ms_s1_chipselect;    // mm_interconnect_0:timer_MS_s1_chipselect -> timer_MS:chipselect
	wire  [15:0] mm_interconnect_0_timer_ms_s1_readdata;      // timer_MS:readdata -> mm_interconnect_0:timer_MS_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_ms_s1_address;       // mm_interconnect_0:timer_MS_s1_address -> timer_MS:address
	wire         mm_interconnect_0_timer_ms_s1_write;         // mm_interconnect_0:timer_MS_s1_write -> timer_MS:write_n
	wire  [15:0] mm_interconnect_0_timer_ms_s1_writedata;     // mm_interconnect_0:timer_MS_s1_writedata -> timer_MS:writedata
	wire         mm_interconnect_0_timer_s_s1_chipselect;     // mm_interconnect_0:timer_S_s1_chipselect -> timer_S:chipselect
	wire  [15:0] mm_interconnect_0_timer_s_s1_readdata;       // timer_S:readdata -> mm_interconnect_0:timer_S_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s_s1_address;        // mm_interconnect_0:timer_S_s1_address -> timer_S:address
	wire         mm_interconnect_0_timer_s_s1_write;          // mm_interconnect_0:timer_S_s1_write -> timer_S:write_n
	wire  [15:0] mm_interconnect_0_timer_s_s1_writedata;      // mm_interconnect_0:timer_S_s1_writedata -> timer_S:writedata
	wire         mm_interconnect_0_button_s1_chipselect;      // mm_interconnect_0:button_s1_chipselect -> button:chipselect
	wire  [31:0] mm_interconnect_0_button_s1_readdata;        // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire   [1:0] mm_interconnect_0_button_s1_address;         // mm_interconnect_0:button_s1_address -> button:address
	wire         mm_interconnect_0_button_s1_write;           // mm_interconnect_0:button_s1_write -> button:write_n
	wire  [31:0] mm_interconnect_0_button_s1_writedata;       // mm_interconnect_0:button_s1_writedata -> button:writedata
	wire         mm_interconnect_0_timer_min_s1_chipselect;   // mm_interconnect_0:timer_min_s1_chipselect -> timer_min:chipselect
	wire  [15:0] mm_interconnect_0_timer_min_s1_readdata;     // timer_min:readdata -> mm_interconnect_0:timer_min_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_min_s1_address;      // mm_interconnect_0:timer_min_s1_address -> timer_min:address
	wire         mm_interconnect_0_timer_min_s1_write;        // mm_interconnect_0:timer_min_s1_write -> timer_min:write_n
	wire  [15:0] mm_interconnect_0_timer_min_s1_writedata;    // mm_interconnect_0:timer_min_s1_writedata -> timer_min:writedata
	wire         mm_interconnect_0_segmentos_5_s1_chipselect; // mm_interconnect_0:segmentos_5_s1_chipselect -> segmentos_5:chipselect
	wire  [31:0] mm_interconnect_0_segmentos_5_s1_readdata;   // segmentos_5:readdata -> mm_interconnect_0:segmentos_5_s1_readdata
	wire   [1:0] mm_interconnect_0_segmentos_5_s1_address;    // mm_interconnect_0:segmentos_5_s1_address -> segmentos_5:address
	wire         mm_interconnect_0_segmentos_5_s1_write;      // mm_interconnect_0:segmentos_5_s1_write -> segmentos_5:write_n
	wire  [31:0] mm_interconnect_0_segmentos_5_s1_writedata;  // mm_interconnect_0:segmentos_5_s1_writedata -> segmentos_5:writedata
	wire         mm_interconnect_0_segmentos_6_s1_chipselect; // mm_interconnect_0:segmentos_6_s1_chipselect -> segmentos_6:chipselect
	wire  [31:0] mm_interconnect_0_segmentos_6_s1_readdata;   // segmentos_6:readdata -> mm_interconnect_0:segmentos_6_s1_readdata
	wire   [1:0] mm_interconnect_0_segmentos_6_s1_address;    // mm_interconnect_0:segmentos_6_s1_address -> segmentos_6:address
	wire         mm_interconnect_0_segmentos_6_s1_write;      // mm_interconnect_0:segmentos_6_s1_write -> segmentos_6:write_n
	wire  [31:0] mm_interconnect_0_segmentos_6_s1_writedata;  // mm_interconnect_0:segmentos_6_s1_writedata -> segmentos_6:writedata
	wire  [31:0] cpu_instruction_master_readdata;             // mm_interconnect_1:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;          // mm_interconnect_1:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [11:0] cpu_instruction_master_address;              // cpu:i_address -> mm_interconnect_1:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                 // cpu:i_read -> mm_interconnect_1:cpu_instruction_master_read
	wire         mm_interconnect_1_rom_s1_chipselect;         // mm_interconnect_1:ROM_s1_chipselect -> ROM:chipselect
	wire  [31:0] mm_interconnect_1_rom_s1_readdata;           // ROM:readdata -> mm_interconnect_1:ROM_s1_readdata
	wire         mm_interconnect_1_rom_s1_debugaccess;        // mm_interconnect_1:ROM_s1_debugaccess -> ROM:debugaccess
	wire   [9:0] mm_interconnect_1_rom_s1_address;            // mm_interconnect_1:ROM_s1_address -> ROM:address
	wire   [3:0] mm_interconnect_1_rom_s1_byteenable;         // mm_interconnect_1:ROM_s1_byteenable -> ROM:byteenable
	wire         mm_interconnect_1_rom_s1_write;              // mm_interconnect_1:ROM_s1_write -> ROM:write
	wire  [31:0] mm_interconnect_1_rom_s1_writedata;          // mm_interconnect_1:ROM_s1_writedata -> ROM:writedata
	wire         mm_interconnect_1_rom_s1_clken;              // mm_interconnect_1:ROM_s1_clken -> ROM:clken
	wire         irq_mapper_receiver0_irq;                    // timer_S:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                    // timer_MS:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                    // button:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                    // timer_min:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                 // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;              // rst_controller:reset_out -> [RAM:reset, ROM:reset, button:reset_n, cpu:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, segmentos_1:reset_n, segmentos_2:reset_n, segmentos_3:reset_n, segmentos_4:reset_n, segmentos_5:reset_n, segmentos_6:reset_n, switchs:reset_n, timer_MS:reset_n, timer_S:reset_n, timer_min:reset_n]
	wire         rst_controller_reset_out_reset_req;          // rst_controller:reset_req -> [RAM:reset_req, ROM:reset_req, rst_translator:reset_req_in]

	platform_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	platform_ROM rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_1_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_1_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_1_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_1_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_1_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_1_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_1_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_1_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	platform_button button (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_s1_readdata),   //                    .readdata
		.in_port    (button_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                //                 irq.irq
	);

	platform_cpu cpu (
		.clk           (clk_clk),                            //                       clk.clk
		.reset_n       (~rst_controller_reset_out_reset),    //                     reset.reset_n
		.d_address     (cpu_data_master_address),            //               data_master.address
		.d_byteenable  (cpu_data_master_byteenable),         //                          .byteenable
		.d_read        (cpu_data_master_read),               //                          .read
		.d_readdata    (cpu_data_master_readdata),           //                          .readdata
		.d_waitrequest (cpu_data_master_waitrequest),        //                          .waitrequest
		.d_write       (cpu_data_master_write),              //                          .write
		.d_writedata   (cpu_data_master_writedata),          //                          .writedata
		.i_address     (cpu_instruction_master_address),     //        instruction_master.address
		.i_read        (cpu_instruction_master_read),        //                          .read
		.i_readdata    (cpu_instruction_master_readdata),    //                          .readdata
		.i_waitrequest (cpu_instruction_master_waitrequest), //                          .waitrequest
		.irq           (cpu_irq_irq),                        //                       irq.irq
		.dummy_ci_port ()                                    // custom_instruction_master.readra
	);

	platform_segmentos_1 segmentos_1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_segmentos_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segmentos_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segmentos_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segmentos_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segmentos_1_s1_readdata),   //                    .readdata
		.out_port   (id7_segmentos_1_external_connection_export)   // external_connection.export
	);

	platform_segmentos_1 segmentos_2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_segmentos_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segmentos_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segmentos_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segmentos_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segmentos_2_s1_readdata),   //                    .readdata
		.out_port   (id7_segmentos_2_external_connection_export)   // external_connection.export
	);

	platform_segmentos_1 segmentos_3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_segmentos_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segmentos_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segmentos_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segmentos_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segmentos_3_s1_readdata),   //                    .readdata
		.out_port   (id7_segmentos_3_external_connection_export)   // external_connection.export
	);

	platform_segmentos_1 segmentos_4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_segmentos_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segmentos_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segmentos_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segmentos_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segmentos_4_s1_readdata),   //                    .readdata
		.out_port   (id7_segmentos_4_external_connection_export)   // external_connection.export
	);

	platform_segmentos_1 segmentos_5 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_segmentos_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segmentos_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segmentos_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segmentos_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segmentos_5_s1_readdata),   //                    .readdata
		.out_port   (segmentos_5_external_connection_export)       // external_connection.export
	);

	platform_segmentos_1 segmentos_6 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_segmentos_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segmentos_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segmentos_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segmentos_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segmentos_6_s1_readdata),   //                    .readdata
		.out_port   (segmentos_6_external_connection_export)       // external_connection.export
	);

	platform_switchs switchs (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_switchs_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switchs_s1_readdata), //                    .readdata
		.in_port  (switchs_external_connection_export)     // external_connection.export
	);

	platform_timer_MS timer_ms (
		.clk        (clk_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_ms_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_ms_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_ms_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_ms_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_ms_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                  //   irq.irq
	);

	platform_timer_S timer_s (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_s_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	platform_timer_min timer_min (
		.clk        (clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_timer_min_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_min_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_min_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_min_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_min_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                   //   irq.irq
	);

	platform_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                         (clk_clk),                                     //                       clk_0_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),              // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address               (cpu_data_master_address),                     //                 cpu_data_master.address
		.cpu_data_master_waitrequest           (cpu_data_master_waitrequest),                 //                                .waitrequest
		.cpu_data_master_byteenable            (cpu_data_master_byteenable),                  //                                .byteenable
		.cpu_data_master_read                  (cpu_data_master_read),                        //                                .read
		.cpu_data_master_readdata              (cpu_data_master_readdata),                    //                                .readdata
		.cpu_data_master_write                 (cpu_data_master_write),                       //                                .write
		.cpu_data_master_writedata             (cpu_data_master_writedata),                   //                                .writedata
		.button_s1_address                     (mm_interconnect_0_button_s1_address),         //                       button_s1.address
		.button_s1_write                       (mm_interconnect_0_button_s1_write),           //                                .write
		.button_s1_readdata                    (mm_interconnect_0_button_s1_readdata),        //                                .readdata
		.button_s1_writedata                   (mm_interconnect_0_button_s1_writedata),       //                                .writedata
		.button_s1_chipselect                  (mm_interconnect_0_button_s1_chipselect),      //                                .chipselect
		.RAM_s1_address                        (mm_interconnect_0_ram_s1_address),            //                          RAM_s1.address
		.RAM_s1_write                          (mm_interconnect_0_ram_s1_write),              //                                .write
		.RAM_s1_readdata                       (mm_interconnect_0_ram_s1_readdata),           //                                .readdata
		.RAM_s1_writedata                      (mm_interconnect_0_ram_s1_writedata),          //                                .writedata
		.RAM_s1_byteenable                     (mm_interconnect_0_ram_s1_byteenable),         //                                .byteenable
		.RAM_s1_chipselect                     (mm_interconnect_0_ram_s1_chipselect),         //                                .chipselect
		.RAM_s1_clken                          (mm_interconnect_0_ram_s1_clken),              //                                .clken
		.segmentos_1_s1_address                (mm_interconnect_0_segmentos_1_s1_address),    //                  segmentos_1_s1.address
		.segmentos_1_s1_write                  (mm_interconnect_0_segmentos_1_s1_write),      //                                .write
		.segmentos_1_s1_readdata               (mm_interconnect_0_segmentos_1_s1_readdata),   //                                .readdata
		.segmentos_1_s1_writedata              (mm_interconnect_0_segmentos_1_s1_writedata),  //                                .writedata
		.segmentos_1_s1_chipselect             (mm_interconnect_0_segmentos_1_s1_chipselect), //                                .chipselect
		.segmentos_2_s1_address                (mm_interconnect_0_segmentos_2_s1_address),    //                  segmentos_2_s1.address
		.segmentos_2_s1_write                  (mm_interconnect_0_segmentos_2_s1_write),      //                                .write
		.segmentos_2_s1_readdata               (mm_interconnect_0_segmentos_2_s1_readdata),   //                                .readdata
		.segmentos_2_s1_writedata              (mm_interconnect_0_segmentos_2_s1_writedata),  //                                .writedata
		.segmentos_2_s1_chipselect             (mm_interconnect_0_segmentos_2_s1_chipselect), //                                .chipselect
		.segmentos_3_s1_address                (mm_interconnect_0_segmentos_3_s1_address),    //                  segmentos_3_s1.address
		.segmentos_3_s1_write                  (mm_interconnect_0_segmentos_3_s1_write),      //                                .write
		.segmentos_3_s1_readdata               (mm_interconnect_0_segmentos_3_s1_readdata),   //                                .readdata
		.segmentos_3_s1_writedata              (mm_interconnect_0_segmentos_3_s1_writedata),  //                                .writedata
		.segmentos_3_s1_chipselect             (mm_interconnect_0_segmentos_3_s1_chipselect), //                                .chipselect
		.segmentos_4_s1_address                (mm_interconnect_0_segmentos_4_s1_address),    //                  segmentos_4_s1.address
		.segmentos_4_s1_write                  (mm_interconnect_0_segmentos_4_s1_write),      //                                .write
		.segmentos_4_s1_readdata               (mm_interconnect_0_segmentos_4_s1_readdata),   //                                .readdata
		.segmentos_4_s1_writedata              (mm_interconnect_0_segmentos_4_s1_writedata),  //                                .writedata
		.segmentos_4_s1_chipselect             (mm_interconnect_0_segmentos_4_s1_chipselect), //                                .chipselect
		.segmentos_5_s1_address                (mm_interconnect_0_segmentos_5_s1_address),    //                  segmentos_5_s1.address
		.segmentos_5_s1_write                  (mm_interconnect_0_segmentos_5_s1_write),      //                                .write
		.segmentos_5_s1_readdata               (mm_interconnect_0_segmentos_5_s1_readdata),   //                                .readdata
		.segmentos_5_s1_writedata              (mm_interconnect_0_segmentos_5_s1_writedata),  //                                .writedata
		.segmentos_5_s1_chipselect             (mm_interconnect_0_segmentos_5_s1_chipselect), //                                .chipselect
		.segmentos_6_s1_address                (mm_interconnect_0_segmentos_6_s1_address),    //                  segmentos_6_s1.address
		.segmentos_6_s1_write                  (mm_interconnect_0_segmentos_6_s1_write),      //                                .write
		.segmentos_6_s1_readdata               (mm_interconnect_0_segmentos_6_s1_readdata),   //                                .readdata
		.segmentos_6_s1_writedata              (mm_interconnect_0_segmentos_6_s1_writedata),  //                                .writedata
		.segmentos_6_s1_chipselect             (mm_interconnect_0_segmentos_6_s1_chipselect), //                                .chipselect
		.switchs_s1_address                    (mm_interconnect_0_switchs_s1_address),        //                      switchs_s1.address
		.switchs_s1_readdata                   (mm_interconnect_0_switchs_s1_readdata),       //                                .readdata
		.timer_min_s1_address                  (mm_interconnect_0_timer_min_s1_address),      //                    timer_min_s1.address
		.timer_min_s1_write                    (mm_interconnect_0_timer_min_s1_write),        //                                .write
		.timer_min_s1_readdata                 (mm_interconnect_0_timer_min_s1_readdata),     //                                .readdata
		.timer_min_s1_writedata                (mm_interconnect_0_timer_min_s1_writedata),    //                                .writedata
		.timer_min_s1_chipselect               (mm_interconnect_0_timer_min_s1_chipselect),   //                                .chipselect
		.timer_MS_s1_address                   (mm_interconnect_0_timer_ms_s1_address),       //                     timer_MS_s1.address
		.timer_MS_s1_write                     (mm_interconnect_0_timer_ms_s1_write),         //                                .write
		.timer_MS_s1_readdata                  (mm_interconnect_0_timer_ms_s1_readdata),      //                                .readdata
		.timer_MS_s1_writedata                 (mm_interconnect_0_timer_ms_s1_writedata),     //                                .writedata
		.timer_MS_s1_chipselect                (mm_interconnect_0_timer_ms_s1_chipselect),    //                                .chipselect
		.timer_S_s1_address                    (mm_interconnect_0_timer_s_s1_address),        //                      timer_S_s1.address
		.timer_S_s1_write                      (mm_interconnect_0_timer_s_s1_write),          //                                .write
		.timer_S_s1_readdata                   (mm_interconnect_0_timer_s_s1_readdata),       //                                .readdata
		.timer_S_s1_writedata                  (mm_interconnect_0_timer_s_s1_writedata),      //                                .writedata
		.timer_S_s1_chipselect                 (mm_interconnect_0_timer_s_s1_chipselect)      //                                .chipselect
	);

	platform_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                         (clk_clk),                              //                       clk_0_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),       // cpu_reset_reset_bridge_in_reset.reset
		.cpu_instruction_master_address        (cpu_instruction_master_address),       //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),   //                                .waitrequest
		.cpu_instruction_master_read           (cpu_instruction_master_read),          //                                .read
		.cpu_instruction_master_readdata       (cpu_instruction_master_readdata),      //                                .readdata
		.ROM_s1_address                        (mm_interconnect_1_rom_s1_address),     //                          ROM_s1.address
		.ROM_s1_write                          (mm_interconnect_1_rom_s1_write),       //                                .write
		.ROM_s1_readdata                       (mm_interconnect_1_rom_s1_readdata),    //                                .readdata
		.ROM_s1_writedata                      (mm_interconnect_1_rom_s1_writedata),   //                                .writedata
		.ROM_s1_byteenable                     (mm_interconnect_1_rom_s1_byteenable),  //                                .byteenable
		.ROM_s1_chipselect                     (mm_interconnect_1_rom_s1_chipselect),  //                                .chipselect
		.ROM_s1_clken                          (mm_interconnect_1_rom_s1_clken),       //                                .clken
		.ROM_s1_debugaccess                    (mm_interconnect_1_rom_s1_debugaccess)  //                                .debugaccess
	);

	platform_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
